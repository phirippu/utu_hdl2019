/home/phil/git/utu_hdl2019/lab_5/lab_5.srcs/sources_1/new/clk_div_4bit.vhd